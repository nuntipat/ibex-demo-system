`ifndef SHUFFLEV_CONSTANT_SV
`define SHUFFLEV_CONSTANT_SV

typedef enum integer {
  RandomSim    = 0,
  RandomTkacik = 1
} shufflev_rng_e;

`endif
